`timescale 1ns / 1ps
module tb();

reg clk, rst, din_rdy, ogot;
reg [31:0] I1, I2;
reg [31:0] i, k; //
wire out_rdy, o_got, gotit, rdy;
wire [31:0] dout;
assign o_got = ogot;
matmult dut(
        .clk(clk),
        .rst(rst),
        .a(I1), 
        .b(I2), 
        .i_ready(din_rdy), 
        .o_got(o_got), 
        .r(dout), 
        .out_ready(out_rdy),
        .gotit(gotit),
        .rdy(rdy));




reg [31:0]din_1[15:0];  // A
reg [31:0]din_2[15:0], save[15:0];  // B
reg [31:0]out[15:0];    // check the result

initial 
begin

   clk <= 1'b0;
   rst <= #10 1'b1;
   rst = #30 1'b0;
   
   i = 32'd0;
  
   din_1[0] = 32'b00111111100000000000000000000000; //1;
   din_2[0] = 32'b00111111100000000000000000000000; //1;
   out[0] = 32'b00111111100000000000000000000000; 
   
   din_1[1] = 32'b00000000000000000000000000000000;//0;
   din_2[1] = 32'b01000000000000000000000000000000; //2;
   out[1] = 32'b01000000000000000000000000000000;
   
   din_1[2] = 32'b00000000000000000000000000000000;//0;
   din_2[2] = 32'b01000000010000000000000000000000;//3;
   out[2] = 32'b01000000010000000000000000000000;
   
   din_1[3] = 32'b00000000000000000000000000000000;//0;
   din_2[3] = 32'b01000000100000000000000000000000;//4
   out[3] = 32'b01000000100000000000000000000000;
   
   din_1[4] = 32'b00000000000000000000000000000000;//0;
   din_2[4] = 32'b00111111100000000000000000000000; //1;
   out[4] = 32'b00111111100000000000000000000000;
   
   din_1[5] = 32'b00111111100000000000000000000000; //1;
   din_2[5] =  32'b01000000000000000000000000000000; //2;
   out[5] = 32'b01000000000000000000000000000000;
   
   din_1[6] = 32'b00000000000000000000000000000000;//0;
   din_2[6] = 32'b01000000010000000000000000000000;//3;
   out[6] = 32'b01000000010000000000000000000000;
   
   din_1[7] = 32'b00000000000000000000000000000000;//0;
   din_2[7] = 32'b01000000100000000000000000000000;//4
   out[7] = 32'b01000000100000000000000000000000;
   
   din_1[8] = 32'b00000000000000000000000000000000;//0;
   din_2[8] = 32'b00111111100000000000000000000000;//1
   out[8] = 32'b00111111100000000000000000000000;
   
   din_1[9] = 32'b00000000000000000000000000000000;//0;
   din_2[9] =  32'b01000000000000000000000000000000; //2;
   out[9] = 32'b01000000000000000000000000000000;
   
   din_1[10] = 32'b00111111100000000000000000000000; //1;
   din_2[10] = 32'b01000000010000000000000000000000;//3;
   out[10] = 32'b01000000010000000000000000000000;
   
   din_1[11] = 32'b00000000000000000000000000000000;//0;
   din_2[11] = 32'b01000000100000000000000000000000;//4
   out[11] = 32'b01000000100000000000000000000000;
   
   din_1[12] = 32'b00000000000000000000000000000000;//0;
   din_2[12] = 32'b00111111100000000000000000000000; //1;
   out[12] = 32'b00111111100000000000000000000000;
   
   din_1[13] = 32'b00000000000000000000000000000000;//0
   din_2[13] =  32'b01000000000000000000000000000000; //2;
   out[13] = 32'b01000000000000000000000000000000;
   
   din_1[14] = 32'b00000000000000000000000000000000;//0;
   din_2[14] = 32'b01000000010000000000000000000000;//3;
   out[14] = 32'b01000000010000000000000000000000;
   
   din_1[15] = 32'b00111111100000000000000000000000;//1
   din_2[15] = 32'b01000000100000000000000000000000;//4
   out[15] = 32'b01000000100000000000000000000000;
   
    /*I1 <= din_1[i];
    I2 <= din_2[i];
    i = i + 1;
    din_rdy <= 1'b1;
    while(gotit != 1'b0)begin end
    din_rdy <= 1'b0;*/
   
   while(i<32'd16)
   begin
        
                ogot <= 1'b1;
                @(posedge rdy) 
                ogot <= 1'b0;               
                I1 <= din_1[i];
                I2 <= din_2[i];
                i=i+1;
                din_rdy <= 1'b1;
                @(posedge gotit) 
                din_rdy <= 1'b0;
            
   end
   
   i = 0;
   ogot <= 1'b1;
   k = 0;
   while(i<32'd16) begin
   
                @(posedge out_rdy);
                ogot <= 1'b0;
                din_rdy <= 1'b1;
                @(posedge gotit)  
                din_rdy <= 1'b0; 
                save[i] <= dout;           
                
                
                if(k == 0)
                    k = k + 1;
                else    
                    i = i+1;
                ogot <= 1'b1;
                
   end
   i = 0;
   while(i<32'd16) begin
        if(save[i]!=out[i])                 
            $display("fail on ",i);
        i = i + 1;
        
   end
end

    always begin 
        #10 clk <= !clk; 
    end

endmodule